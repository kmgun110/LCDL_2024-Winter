//This is for the 4:2 priority encoder module.

module four_to_two_priority_encoder_dataflow_module (a, b, c, d, out0, out1);
	input a, b, c, d;

	output out0, out1;

	assign out0 = d || (b && !c);
	assign out1 = c || d;

endmodule


